//
// University of Utah, Computer Design Laboratory ECE 3710, CompactRISC16
//
// Create Date: 10/08/2021
// Module Name: cr16
// Description: The CompactRISC16 (CR16) processor with an integrated FSM and instruction decoder
// along with an instantiated datapath, ALU, and program counter.
// Authors: Jacob Peterson, Brady Hartog, Isabella Gilman, Nate Hansen
//

module cr16 ();

// TODO implement CR16 decoder and FSM, instantiate other modules
// This should not instantiate BRAM, but rather have port interfaces for it
// so that a memory mapping module (for virtual memory addressing or mapping certain addresses to
// a peripheral register/interface) can be used outside of this project.

endmodule
