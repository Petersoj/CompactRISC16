//
// University of Utah, Computer Design Laboratory ECE 3710, CompactRISC16
//
// Create Date: 10/7/2021
// Module Name: pc
// Description: Program counter to drive the FSM of the CR16 ALU. 
// Authors: Jacob Peterson, Brady Hartog, Isabella Gilman, Nate Hansen
//