//
// University of Utah, Computer Design Laboratory ECE 3710, CompactRISC16
//
// Create Date: 10/7/2021
// Module Name: decoder
// Description: 
// Authors: Jacob Peterson, Brady Hartog, Isabella Gilman, Nate Hansen
//

